// Drake Gonzales
// drgonzales@g.hmc.edu
// This Module holds the mixcol module
// 11/03/25

module mixcolumn(input  logic [31:0] a,
                 input  logic  alarm,
                 output logic [31:0] y);
                      

    logic [7:0] a0, a1, a2, a3, y0, y1, y2, y3, t0, t1, t2, t3, tmp;
    logic [31:0] mix_result;
        assign {a0, a1, a2, a3} = a;
        assign tmp = a0 ^ a1 ^ a2 ^ a3;
    
        galoismult gm0(a0^a1, t0);
        galoismult gm1(a1^a2, t1);
        galoismult gm2(a2^a3, t2);
        galoismult gm3(a3^a0, t3);
        
        assign y0 = a0 ^ tmp ^ t0;
        assign y1 = a1 ^ tmp ^ t1;
        assign y2 = a2 ^ tmp ^ t2;
        assign y3 = a3 ^ tmp ^ t3;
        assign mix_result = {y0, y1, y2, y3}; 

        assign y = (alarm == 1'b1) ? a : mix_result;
        

endmodule